library verilog;
use verilog.vl_types.all;
entity lfsr5b_tb is
end lfsr5b_tb;
