library verilog;
use verilog.vl_types.all;
entity bist_tb is
end bist_tb;
