library verilog;
use verilog.vl_types.all;
entity ex2_tb is
end ex2_tb;
