library verilog;
use verilog.vl_types.all;
entity sisr4b_tb is
end sisr4b_tb;
