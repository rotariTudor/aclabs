library verilog;
use verilog.vl_types.all;
entity fdivby5_tb is
end fdivby5_tb;
