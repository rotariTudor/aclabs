library verilog;
use verilog.vl_types.all;
entity fsm_1011_tb is
end fsm_1011_tb;
