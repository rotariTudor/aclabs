library verilog;
use verilog.vl_types.all;
entity lfsr_tb is
end lfsr_tb;
