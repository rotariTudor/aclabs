library verilog;
use verilog.vl_types.all;
entity check_tb is
end check_tb;
