library verilog;
use verilog.vl_types.all;
entity ex3_tb is
end ex3_tb;
