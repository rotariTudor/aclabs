library verilog;
use verilog.vl_types.all;
entity tb_comp_3b is
end tb_comp_3b;
