library verilog;
use verilog.vl_types.all;
entity regfl_4x8_tb is
end regfl_4x8_tb;
