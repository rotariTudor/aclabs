library verilog;
use verilog.vl_types.all;
entity r4b_tb is
end r4b_tb;
