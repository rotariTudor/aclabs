library verilog;
use verilog.vl_types.all;
entity cmp4b_tb is
end cmp4b_tb;
