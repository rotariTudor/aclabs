library verilog;
use verilog.vl_types.all;
entity hotfsm_tb is
end hotfsm_tb;
