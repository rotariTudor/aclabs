library verilog;
use verilog.vl_types.all;
entity ex1a_tb is
end ex1a_tb;
