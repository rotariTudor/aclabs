library verilog;
use verilog.vl_types.all;
entity div3_tb is
end div3_tb;
