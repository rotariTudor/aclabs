library verilog;
use verilog.vl_types.all;
entity cnt1s_tb is
end cnt1s_tb;
