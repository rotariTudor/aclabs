module lfsr