library verilog;
use verilog.vl_types.all;
entity fdivby3_tb is
end fdivby3_tb;
