library verilog;
use verilog.vl_types.all;
entity sadd_tb is
end sadd_tb;
