library verilog;
use verilog.vl_types.all;
entity karnaugh_tb is
end karnaugh_tb;
