library verilog;
use verilog.vl_types.all;
entity dec2x4_tb is
end dec2x4_tb;
