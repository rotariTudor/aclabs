library verilog;
use verilog.vl_types.all;
entity fac_tb is
end fac_tb;
