library verilog;
use verilog.vl_types.all;
entity mlopadd_tb is
end mlopadd_tb;
