library verilog;
use verilog.vl_types.all;
entity ex1a is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        f1              : out    vl_logic
    );
end ex1a;
