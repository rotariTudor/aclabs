library verilog;
use verilog.vl_types.all;
entity add2b_tb is
end add2b_tb;
