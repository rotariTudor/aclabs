library verilog;
use verilog.vl_types.all;
entity ex4_tb is
end ex4_tb;
